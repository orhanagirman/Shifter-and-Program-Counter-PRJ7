----------------------------------------------------------------------------------
-- Company: 
-- Engineer: 
-- 
-- Create Date:    14:07:12 08/07/2020 
-- Design Name: 
-- Module Name:    fulladder - Behavioral 
-- Project Name: 
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity fulladder is
    Port ( a : in  STD_LOGIC;
           b : in   STD_LOGIC;
           cin : in  STD_LOGIC;
			  cout : out STD_LOGIC;
           s : out  STD_LOGIC);
end fulladder;

architecture Behavioral of fulladder is

signal wire1 : STD_LOGIC;
signal wire2 : STD_LOGIC;
signal wire3 : STD_LOGIC;

begin
     
	  wire1 <= a xor b ;
	  wire2 <= a and b ;
	  s <= wire1 xor cin ;
	  wire3 <= wire1 and cin ;
	  cout <= wire2 or wire3 ;

			
end Behavioral;

